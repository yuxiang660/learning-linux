module tb;

initial
   begin
      $display("Hello World!");
   end

endmodule
